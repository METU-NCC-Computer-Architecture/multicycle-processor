library verilog;
use verilog.vl_types.all;
entity SHIFTREG8_vlg_vec_tst is
end SHIFTREG8_vlg_vec_tst;
