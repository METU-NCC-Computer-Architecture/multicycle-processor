library verilog;
use verilog.vl_types.all;
entity SHIFTREGS_vlg_vec_tst is
end SHIFTREGS_vlg_vec_tst;
