library verilog;
use verilog.vl_types.all;
entity MUX2TO1_vlg_vec_tst is
end MUX2TO1_vlg_vec_tst;
