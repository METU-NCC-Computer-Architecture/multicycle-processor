library verilog;
use verilog.vl_types.all;
entity ap_function_vlg_vec_tst is
end ap_function_vlg_vec_tst;
