library verilog;
use verilog.vl_types.all;
entity deneme_vlg_vec_tst is
end deneme_vlg_vec_tst;
