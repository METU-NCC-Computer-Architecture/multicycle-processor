library verilog;
use verilog.vl_types.all;
entity DFF8_vlg_vec_tst is
end DFF8_vlg_vec_tst;
