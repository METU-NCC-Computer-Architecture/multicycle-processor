library verilog;
use verilog.vl_types.all;
entity SIGNEXT6T08_vlg_vec_tst is
end SIGNEXT6T08_vlg_vec_tst;
