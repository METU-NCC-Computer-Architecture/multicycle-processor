library verilog;
use verilog.vl_types.all;
entity Datapath is
    port(
        altera_reserved_tms: in     vl_logic;
        altera_reserved_tck: in     vl_logic;
        altera_reserved_tdi: in     vl_logic;
        altera_reserved_tdo: out    vl_logic;
        Qm1             : out    vl_logic;
        RST             : in     vl_logic;
        LDQ             : in     vl_logic;
        CLK             : in     vl_logic;
        LDA             : in     vl_logic;
        A               : out    vl_logic_vector(7 downto 0);
        SR_SEL          : in     vl_logic;
        MULT_SEL        : in     vl_logic;
        Cin             : in     vl_logic;
        PC_EN           : in     vl_logic;
        INST_MEM_OUT    : in     vl_logic_vector(15 downto 0);
        PC_MUX_SEL      : in     vl_logic_vector(1 downto 0);
        RF_EN           : in     vl_logic;
        INS_TYPE_MUX_SEL: in     vl_logic;
        PLUS1_SEL       : in     vl_logic;
        DATA_MEM_OUT    : in     vl_logic_vector(15 downto 0);
        D_SEL           : in     vl_logic_vector(1 downto 0);
        A_SEL           : in     vl_logic_vector(1 downto 0);
        OAP             : in     vl_logic_vector(2 downto 0);
        B_SEL           : in     vl_logic_vector(1 downto 0);
        Product         : out    vl_logic_vector(15 downto 0);
        MULT_EN         : in     vl_logic;
        SR              : in     vl_logic;
        SL              : in     vl_logic;
        CO              : out    vl_logic;
        OVF             : out    vl_logic;
        Z               : out    vl_logic;
        N               : out    vl_logic;
        ALUOUT          : out    vl_logic_vector(7 downto 0);
        OPCODE          : out    vl_logic_vector(3 downto 0);
        OUT_Q           : out    vl_logic_vector(7 downto 0);
        READ_DATA_A     : out    vl_logic_vector(7 downto 0);
        READ_DATA_B     : out    vl_logic_vector(7 downto 0);
        RF_OUT_A        : out    vl_logic_vector(7 downto 0);
        RF_OUT_B        : out    vl_logic_vector(7 downto 0);
        RF_R_ADDR_B     : out    vl_logic_vector(2 downto 0);
        RF_W_ADDR       : out    vl_logic_vector(2 downto 0);
        RF_W_DATA       : out    vl_logic_vector(7 downto 0);
        WB_SEL          : in     vl_logic;
        UL_SEL          : in     vl_logic
    );
end Datapath;
