library verilog;
use verilog.vl_types.all;
entity RegisterFile8x8_vlg_vec_tst is
end RegisterFile8x8_vlg_vec_tst;
