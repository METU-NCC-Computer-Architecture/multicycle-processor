library verilog;
use verilog.vl_types.all;
entity ROUTER_vlg_vec_tst is
end ROUTER_vlg_vec_tst;
