library verilog;
use verilog.vl_types.all;
entity MUX4TO1_vlg_vec_tst is
end MUX4TO1_vlg_vec_tst;
