library verilog;
use verilog.vl_types.all;
entity simple_divider_vlg_vec_tst is
end simple_divider_vlg_vec_tst;
